package agent_pkg;
  import uvm_pkg::*;
  `include "packet.sv"
  `include "packet2.sv"
  `include "monitor.sv"
  `include "driver.sv"
  `include "agent.sv"
  `include "output_packet.sv"
  `include "output_monitor.sv"
  `include "output_agent.sv"

endpackage
